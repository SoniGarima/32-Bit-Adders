`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.10.2019 22:15:23
// Design Name: 
// Module Name: cla32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cla32(
    input [31:0] A,
    input [31:0] B,
    input Cin,
    output [32:0] Sum,
    output Cout
    );
    wire [31:0] P,G,C;
    assign P=A^B;
    assign G=A&B;
 assign C[0]=Cin;
 assign C[1]=(G[0]|P[0]&Cin);
assign C[2]=(G[1]|P[1]&(G[0]|P[0]&Cin));
assign C[3]=(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)));
assign C[4]=(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))));
assign C[5]=(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))));
assign C[6]=(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))));
assign C[7]=(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))));
assign C[8]=(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))));
assign C[9]=(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))));
assign C[10]=(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))));
assign C[11]=(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))));
assign C[12]=(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))));
assign C[13]=(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))));
assign C[14]=(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))));
assign C[15]=(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))));
assign C[16]=(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))));
assign C[17]=(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))));
assign C[18]=(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))));
assign C[19]=(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))));
assign C[20]=(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))));
assign C[21]=(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))));
assign C[22]=(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))));
assign C[23]=(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))))));
assign C[24]=(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))))));
assign C[25]=(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))))))));
assign C[26]=(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))))))));
assign C[27]=(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))))))))));
assign C[28]=(G[27]|P[27]&(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))))))))));
assign C[29]=(G[28]|P[28]&(G[27]|P[27]&(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))))))))))));
assign C[30]=(G[29]|P[29]&(G[28]|P[28]&(G[27]|P[27]&(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))))))))))));
assign C[31]=(G[30]|P[30]&(G[29]|P[29]&(G[28]|P[28]&(G[27]|P[27]&(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin)))))))))))))))))))))))))))))));
assign Cout=(G[31]|P[31]&(G[30]|P[30]&(G[29]|P[29]&(G[28]|P[28]&(G[27]|P[27]&(G[26]|P[26]&(G[25]|P[25]&(G[24]|P[24]&(G[23]|P[23]&(G[22]|P[22]&(G[21]|P[21]&(G[20]|P[20]&(G[19]|P[19]&(G[18]|P[18]&(G[17]|P[17]&(G[16]|P[16]&(G[15]|P[15]&(G[14]|P[14]&(G[13]|P[13]&(G[12]|P[12]&(G[11]|P[11]&(G[10]|P[10]&(G[9]|P[9]&(G[8]|P[8]&(G[7]|P[7]&(G[6]|P[6]&(G[5]|P[5]&(G[4]|P[4]&(G[3]|P[3]&(G[2]|P[2]&(G[1]|P[1]&(G[0]|P[0]&Cin))))))))))))))))))))))))))))))));
assign Sum=C^A^B;
assign Sum[32]=Cout;
endmodule
